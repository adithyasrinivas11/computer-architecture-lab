`include "mux2.v"

module barelshift (s,inp,outp);
	input [3:0]s;
	wire s0,s1,s2,s3,s4;
	input [15:0] inp;
	output [15:0] outp;
	wire [15:0] w1,w2,w3,w4;

assign s0=s[0];
assign s1=s[1];
assign s2=s[2];
assign s3=s[3];

mux_2_1_1 m1(s0,1'b0,inp[0],w1[0]);
mux_2_1_1 m11(s0,inp[0],inp[1],w1[1]);
mux_2_1_1 m12(s0,inp[1],inp[2],w1[2]);
mux_2_1_1 m13(s0,inp[2],inp[3],w1[3]);
mux_2_1_1 m14(s0,inp[3],inp[4],w1[4]);
mux_2_1_1 m15(s0,inp[4],inp[5],w1[5]);
mux_2_1_1 m16(s0,inp[5],inp[6],w1[6]);
mux_2_1_1 m17(s0,inp[6],inp[7],w1[7]);
mux_2_1_1 m18(s0,inp[7],inp[8],w1[8]);
mux_2_1_1 m19(s0,inp[8],inp[9],w1[9]);
mux_2_1_1 m191(s0,inp[9],inp[10],w1[10]);
mux_2_1_1 m162(s0,inp[10],inp[11],w1[11]);
mux_2_1_1 m1732(s0,inp[11],inp[12],w1[12]);
mux_2_1_1 m1813(s0,inp[12],inp[13],w1[13]);
mux_2_1_1 m1913(s0,inp[13],inp[14],w1[14]);
mux_2_1_1 m1912(s0,inp[14],inp[15],w1[15]);


mux_2_1_1 m20(s1,1'b0,w1[0],w2[0]);
mux_2_1_1 m21(s1,1'b0,w1[1],w2[1]);
mux_2_1_1 m22(s1,w1[0],w1[2],w2[2]);
mux_2_1_1 m23(s1,w1[1],w1[3],w2[3]);
mux_2_1_1 m24(s1,w1[2],w1[4],w2[4]);
mux_2_1_1 m25(s1,w1[3],w1[5],w2[5]);
mux_2_1_1 m26(s1,w1[4],w1[6],w2[6]);
mux_2_1_1 m27(s1,w1[5],w1[7],w2[7]);
mux_2_1_1 m28(s1,w1[6],w1[8],w2[8]);
mux_2_1_1 m29(s1,w1[7],w1[9],w2[9]);
mux_2_1_1 m291(s1,w1[8],w1[10],w2[10]);
mux_2_1_1 m230(s1,w1[9],w1[11],w2[11]);
mux_2_1_1 m240(s1,w1[10],w1[12],w2[12]);
mux_2_1_1 m250(s1,w1[11],w1[13],w2[13]);
mux_2_1_1 m260(s1,w1[12],w1[14],w2[14]);
mux_2_1_1 m270(s1,w1[13],w1[15],w2[15]);


mux_2_1_1 m40(s2,1'b0,w2[0],w3[0]);
mux_2_1_1 m41(s2,1'b0,w2[1],w3[1]);
mux_2_1_1 m42(s2,1'b0,w2[2],w3[2]);
mux_2_1_1 m43(s2,1'b0,w2[3],w3[3]);
mux_2_1_1 m44(s2,w2[0],w2[4],w3[4]);
mux_2_1_1 m45(s2,w2[1],w2[5],w3[5]);
mux_2_1_1 m46(s2,w2[2],w2[6],w3[6]);
mux_2_1_1 m47(s2,w2[3],w2[7],w3[7]);
mux_2_1_1 m48(s2,w2[4],w2[8],w3[8]);
mux_2_1_1 m49(s2,w2[5],w2[9],w3[9]);
mux_2_1_1 m491(s2,w2[6],w2[10],w3[10]);
mux_2_1_1 m441(s2,w2[7],w2[11],w3[11]);
mux_2_1_1 m451(s2,w2[8],w2[12],w3[12]);
mux_2_1_1 m461(s2,w2[9],w2[13],w3[13]);
mux_2_1_1 m471(s2,w2[10],w2[14],w3[14]);
mux_2_1_1 m481(s2,w2[11],w2[15],w3[15]);



mux_2_1_1 m80(s3,1'b0,w3[0],w4[0]);
mux_2_1_1 m81(s3,1'b0,w3[1],w4[1]);
mux_2_1_1 m82(s3,1'b0,w3[2],w4[2]);
mux_2_1_1 m83(s3,1'b0,w3[3],w4[3]);
mux_2_1_1 m84(s3,1'b0,w3[4],w4[4]);
mux_2_1_1 m85(s3,1'b0,w3[5],w4[5]);
mux_2_1_1 m86(s3,1'b0,w3[6],w4[6]);
mux_2_1_1 m87(s3,1'b0,w3[7],w4[7]);
mux_2_1_1 m88(s3,w3[0],w3[8],w4[8]);
mux_2_1_1 m89(s3,w3[1],w3[9],w4[9]);
mux_2_1_1 m891(s3,w3[2],w3[10],w4[10]);
mux_2_1_1 m881(s3,w3[3],w3[11],w4[11]);
mux_2_1_1 m892(s3,w3[4],w3[12],w4[12]);
mux_2_1_1 m8921(s3,w3[5],w3[13],w4[13]);
mux_2_1_1 m882(s3,w3[6],w3[14],w4[14]);
mux_2_1_1 m893(s3,w3[7],w3[15],w4[15]);


assign outp[15:0]=w4[15:0];



endmodule
