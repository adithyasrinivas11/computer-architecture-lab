`include "2x1mux.v"

module bar_shif(s,i,op);

input [3:0]s;
input [15:0]i;

output [15:0]op;

wire [15:0]w1,w2,w3,w4;

mux21 m1(i[0],i[1],s[0],w1[0]); 					//s =1 then i1 is choosen
mux21 m2(i[1],i[2],s[0],w1[1]);
mux21 m3(i[2],i[3],s[0],w1[2]);
mux21 m4(i[3],i[4],s[0],w1[3]);
mux21 m5(i[4],i[5],s[0],w1[4]);
mux21 m6(i[5],i[6],s[0],w1[5]);
mux21 m7(i[6],i[7],s[0],w1[6]);
mux21 m8(i[7],i[8],s[0],w1[7]);
mux21 m9(i[8],i[9],s[0],w1[8]);
mux21 m01(i[9],i[10],s[0],w1[9]);
mux21 m02(i[10],i[11],s[0],w1[10]);
mux21 m03(i[11],i[12],s[0],w1[11]);
mux21 m04(i[12],i[13],s[0],w1[12]);
mux21 m05(i[13],i[14],s[0],w1[13]);
mux21 m06(i[14],i[15],s[0],w1[14]);
mux21 m011(i[15],1'b0,s[0],w1[15]);

mux21 m11(w1[0],w1[2],s[1],w2[0]);
mux21 m12(w1[1],w1[3],s[1],w2[1]);
mux21 m13(w1[2],w1[4],s[1],w2[2]);
mux21 m14(w1[3],w1[5],s[1],w2[3]);
mux21 m15(w1[4],w1[6],s[1],w2[4]);
mux21 m16(w1[5],w1[7],s[1],w2[5]);
mux21 m17(w1[6],w1[8],s[1],w2[6]);
mux21 m18(w1[7],w1[9],s[1],w2[7]);
mux21 m19(w1[8],w1[10],s[1],w2[8]);
mux21 m111(w1[9],w1[11],s[1],w2[9]);
mux21 m121(w1[10],w1[12],s[1],w2[10]);
mux21 m131(w1[11],w1[13],s[1],w2[11]);
mux21 m141(w1[12],w1[14],s[1],w2[12]);
mux21 m151(w1[13],w1[15],s[1],w2[13]);
mux21 m101(w1[14],1'b0,s[1],w2[14]);
mux21 m1011(w1[15],1'b0,s[1],w2[15]);

mux21 m21(w2[0],w2[4],s[2],w3[0]);
mux21 m22(w2[1],w2[5],s[2],w3[1]);
mux21 m23(w2[2],w2[6],s[2],w3[2]);
mux21 m24(w2[3],w2[7],s[2],w3[3]);
mux21 m25(w2[4],w2[8],s[2],w3[4]);
mux21 m26(w2[5],w2[9],s[2],w3[5]);
mux21 m27(w2[6],w2[10],s[2],w3[6]);
mux21 m211(w2[7],w2[11],s[2],w3[7]);
mux21 m221(w2[8],w2[12],s[2],w3[8]);
mux21 m231(w2[9],w2[13],s[2],w3[9]);
mux21 m241(w2[10],w2[14],s[2],w3[10]);
mux21 m251(w2[11],w2[15],s[2],w3[11]);
mux21 m281(w2[12],1'b0,s[2],w3[12]);
mux21 m291(w2[13],1'b0,s[2],w3[13]);
mux21 m201(w2[14],1'b0,s[2],w3[14]);
mux21 m2011(w2[15],1'b0,s[2],w3[15]);

//////////////////////////////////////////////////////////////////////

mux21 m31(w3[0],w3[8],s[3],w4[0]);
mux21 m32(w3[1],w3[9],s[3],w4[1]);
mux21 m33(w3[2],w3[10],s[3],w4[2]);
mux21 m311(w3[3],w3[11],s[3],w4[3]);
mux21 m321(w3[4],w3[12],s[3],w4[4]);
mux21 m331(w3[5],w3[13],s[3],w4[5]);
mux21 m312(w3[6],w3[14],s[3],w4[6]);
mux21 m3121(w3[7],w3[15],s[3],w4[7]);
mux21 m342(w3[8],1'b0,s[3],w4[8]);
mux21 m3523(w3[9],1'b0,s[3],w4[9]);
mux21 m3613(w3[10],1'b0,s[3],w4[10]);
mux21 m3731(w3[11],1'b0,s[3],w4[11]);
mux21 m383(w3[12],1'b0,s[3],w4[12]);
mux21 m394(w3[13],1'b0,s[3],w4[13]);
mux21 m3055(w3[14],1'b0,s[3],w4[14]);
mux21 m311112(w3[15],1'b0,s[3],w4[15]);

assign op[15:0]=w4[15:0];


endmodule
